// -------------------- define timescale -----------------------
`timescale 1ns/1ps

module mux_control_tb();

// -------------------- define parameters -----------------------
parameter NUMSTAGES = 5;
parameter NUMSAMPLES = 32;
parameter WORDSIZE = 16;
parameter WL=16, IWL=5, FWL=10;

// -------------------- create inputs and oututs -----------------------
reg [NUMSTAGES-3:0] counter_r;
reg [2:0] stage_num_r;
wire m0_s, m2_s, m3_s;
wire [1:0] m1_s;

// -------------------- testbench variables -----------------------
reg clk;

// -------------------- module being tested -----------------------
mux_control #(.NUMSTAGES(NUMSTAGES)) m0(
	counter_r,
	stage_num_r,
	m0_s, m1_s, m2_s, m3_s	
);

// -------------------- initialize -----------------------
initial
begin
	clk <= 0;
	counter_r <= 0;
	stage_num_r <= 0;
end

// -------------------- clock generation -----------------------
always @(*)
begin
	clk <= #0.05~clk;
end

// -------------------- testing -----------------------
always @(posedge clk)
begin
	if(stage_num_r < 3'b101)
	begin
		if(counter_r == {NUMSTAGES-2{1'b1}})
		begin
			stage_num_r = stage_num_r + 1;
			counter_r <= 0;
		end else 
			counter_r <= counter_r + 1;
	end
end

endmodule
